module segments_lut(input [4:0] score, output [13:0] segments);
    reg[13:0] seg;
    assign segments = seg;

    always @(score) begin
        case(score)
            5'd0  : seg = 14'b00000000111111;
            5'd1  : seg = 14'b00000000000011;
            5'd2  : seg = 14'b00000001101101;
            5'd3  : seg = 14'b00000001100111;
            5'd4  : seg = 14'b00000001010011;
            5'd5  : seg = 14'b00000001110110;
            5'd6  : seg = 14'b00000001111110;
            5'd7  : seg = 14'b00000000100011;
            5'd8  : seg = 14'b00000001111111;
            5'd9  : seg = 14'b00000001110111;
            5'd10 : seg = 14'b00000110111111;
            5'd11 : seg = 14'b00000110000011;
            5'd12 : seg = 14'b00000111101101;
            5'd13 : seg = 14'b00000111100111;
            5'd14 : seg = 14'b00000111010011;
            5'd15 : seg = 14'b00000111110110;
            5'd16 : seg = 14'b00000111111110;
            5'd17 : seg = 14'b00000110100011;
            5'd18 : seg = 14'b00000111111111;
            5'd19 : seg = 14'b00000111110111;
            5'd20 : seg = 14'b11011010111111;
            5'd21 : seg = 14'b11011010000011;
            5'd22 : seg = 14'b11011011101101;
            5'd23 : seg = 14'b11011011100111;
            5'd24 : seg = 14'b11011011010011;
            5'd25 : seg = 14'b11011011110110;
            5'd26 : seg = 14'b11011011111110;
            5'd27 : seg = 14'b11011010100011;
            5'd28 : seg = 14'b11011011111111;
            5'd29 : seg = 14'b11011011110111;
            5'd30 : seg = 14'b11001110111111;
            5'd31 : seg = 14'b11001110000011;

            default: seg = 7'b00000001111000;
        endcase
    end
endmodule